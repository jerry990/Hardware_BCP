`define Adus  2
`define DATA_SIZE 18
`define ADDR_SIZE 12